//******************************************************************************
// File name        : StrobeGen.v
// Module name      : StrobeGen
// Company          : Radware
// Project name     : ODS-MR
// Card name        : Yarkon
// Designer         : Iris  Bener Sharoni
// Creation Date    : 15.10.2010
// Status           : Under design
// Last modified by : Carlos Chen
// Last modified    : 07.10.2015
// Version          : 1.0
// Description      : Generates cyclic strobe signals
// Hierarchy Up     : ODS_MR
// Hierarchy Down   : -
// Card Release     : 1.0
//******************************************************************************

//------------------------------------------------------------------------------
// Macro define or include file
//------------------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Module declaration
//------------------------------------------------------------------------------
module StrobeGen (
    ResetN,         // In,
    LpcClock,       // In, 33 MHz Lpc (Altera Clock)
    SlowClock,      // In, Oscillator Clock 32,768 Hz
    Strobe1s,       // Out, Single SlowClock Pulse @ 1 s
    Strobe488us,    // Out, Single SlowClock Pulse @ 488 us
    Strobe1ms,      // Out, Single SlowClock Pulse @ 1 ms
    Strobe16ms,     // Out, Single SlowClock Pulse @ 16 ms
    Strobe125ms,    // Out, Single SlowClock Pulse @ 125 ms
    Strobe125msec,  // Out, Single LpcClock  Pulse @ 125 ms
    Counter         // Out, 15 bit Free run Counter on Slow Clock
);

//------------------------------------------------------------------------------
// Parameter declaration
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// User defined parameter
//--------------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Standard parameter
//--------------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Local parameter
//--------------------------------------------------------------------------
// time delay, flip-flop output assignment delay for simulation waveform trace
localparam TD = 1;

//------------------------------------------------------------------------------
// Variable declaration
//------------------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Input/Output declaration
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// Input declaration
//--------------------------------------------------------------------------
input           ResetN;
input           LpcClock;
input           SlowClock;

//--------------------------------------------------------------------------
// Output declaration
//--------------------------------------------------------------------------
output          Strobe1s;
output          Strobe1ms;
output          Strobe16ms;
output          Strobe125ms;
output          Strobe125msec;
output          Strobe488us;
output  [14:0]  Counter;

//------------------------------------------------------------------------------
// Signal declaration
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// Wire declaration
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Combinational, module connection
//----------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Reg declaration
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Combinational
//----------------------------------------------------------------------
//------------------------------------------------------------------
// Output
//------------------------------------------------------------------
// None

//------------------------------------------------------------------
// Internal signal
//------------------------------------------------------------------
// None

//------------------------------------------------------------------
// FSM
//------------------------------------------------------------------
// None

//----------------------------------------------------------------------
// Sequential
//----------------------------------------------------------------------
//------------------------------------------------------------------
// Output
//------------------------------------------------------------------
reg             Strobe1s;
reg             Strobe1ms;
reg             Strobe16ms;
reg             Strobe125ms;
reg             Strobe488us;
reg     [14:0]  Counter;

//------------------------------------------------------------------
// Internal signal
//------------------------------------------------------------------
reg     [1:0]   StrobeEdge;
reg             Strobe125msec;

//------------------------------------------------------------------
// FSM
//------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Task/Function description and included task/function description
//------------------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Main code
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// Combinational circuit
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Output
//----------------------------------------------------------------------
// None

//----------------------------------------------------------------------
// Internal signal
//----------------------------------------------------------------------
// None

//----------------------------------------------------------------------
// FSM
//----------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Sequential circuit
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Output
//----------------------------------------------------------------------
always @ (posedge SlowClock or negedge ResetN) begin
  if (!ResetN) begin
      Strobe1s <= #TD 1'b0;
      Strobe1ms <= #TD 1'b0;
      Strobe16ms <= #TD 1'b0;
      Strobe125ms <= #TD 1'b0;
      Strobe488us <= #TD 1'b0;
      Counter <= #TD 15'd0;
  end else begin
      Strobe1s <= #TD (Counter == 15'h5);
      Strobe1ms <= #TD (Counter[4:0] == 5'h5);
      Strobe16ms <= #TD (Counter[8:0] == 9'h5);
      Strobe125ms <= #TD (Counter[11:0] == 12'h5);
      Strobe488us <= #TD (Counter[3:0] == 4'h5);
      Counter <= #TD Counter + 15'd1;
  end
end

always @ (posedge LpcClock or negedge ResetN) begin
  if (!ResetN)
      Strobe125msec <= #TD 0;
  else
      Strobe125msec <= #TD (StrobeEdge == 2'h1);
end

//----------------------------------------------------------------------
// Internal signal
//----------------------------------------------------------------------
always @ (posedge LpcClock or negedge ResetN) begin
  if (!ResetN)
      StrobeEdge <= #TD 2'b00;
  else
      StrobeEdge <= #TD {StrobeEdge[0], Strobe125ms};
end

//----------------------------------------------------------------------
// FSM
//----------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Module instantiation
//--------------------------------------------------------------------------
// None

endmodule
