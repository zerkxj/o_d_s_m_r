//******************************************************************************
// File name        : PwrBtnControl.v
// Module name      : PwrBtnControl
// Description      : This module control Power Btuuon timing
// Hierarchy Up     : ODS_MR
// Hierarchy Down   : ---
//******************************************************************************

//------------------------------------------------------------------------------
// Macro define or include file
//------------------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Module declaration
//------------------------------------------------------------------------------
module  PwrBtnControl (
    InitResetN,         // In,
    Strobe125ms,        // In,
    PWR_BTN_IN_N,       // In,
    PWRGD_PS_PWROK_3V3, // In,
    FM_PS_EN,           // In,
    PowerEvtState,      // In,
    PowerButtonOut_ox,  // In,
    PowerbuttonEvtOut,  // In,
    RstBiosFlg,         // Out,
    FM_SYS_SIO_PWRBTN_N // Out
);


//------------------------------------------------------------------------------
// Parameter declaration
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// User defined parameter
//--------------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Standard parameter
//--------------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Local parameter
//--------------------------------------------------------------------------
// time delay, flip-flop output assignment delay for simulation waveform trace
localparam TD = 1;

//------------------------------------------------------------------------------
// Variable declaration
//------------------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Input/Output declaration
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// Input declaration
//--------------------------------------------------------------------------
input           InitResetN;
input           Strobe125ms;
input           PWR_BTN_IN_N;
input           PWRGD_PS_PWROK_3V3;
input           FM_PS_EN;
input   [3:0]   PowerEvtState;
input           PowerButtonOut_ox;  // From MR_Bsp.ButtonControl.Button::StrobeOut ( in ButtonControl.v file )
input           PowerbuttonEvtOut;  // From PwrEvent

//--------------------------------------------------------------------------
// Output declaration
//--------------------------------------------------------------------------
output          RstBiosFlg; // To MR_Bsp.BiosControl
output          FM_SYS_SIO_PWRBTN_N; // Output to SIO

//------------------------------------------------------------------------------
// Signal declaration
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// Wire declaration
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Combinational, module connection
//----------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Reg declaration
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Combinational
//----------------------------------------------------------------------
//------------------------------------------------------------------
// Output
//------------------------------------------------------------------
// None

//------------------------------------------------------------------
// Internal signal
//------------------------------------------------------------------
// None

//------------------------------------------------------------------
// FSM
//------------------------------------------------------------------
// None

//----------------------------------------------------------------------
// Sequential
//----------------------------------------------------------------------
//------------------------------------------------------------------
// Output
//------------------------------------------------------------------
// None

//------------------------------------------------------------------
// Internal signal
//------------------------------------------------------------------
reg     [9:0]   PowerButtonInBuf;

//------------------------------------------------------------------
// FSM
//------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Task/Function description and included task/function description
//------------------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Main code
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// Combinational circuit
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Output
//----------------------------------------------------------------------
assign RstBiosFlg = (PWRGD_PS_PWROK_3V3) ? 1'b0 :
                        ((PowerEvtState == `Event_PowerStandBy) && (~PWR_BTN_IN_N)) ? 1'b1 :
                            ((~PowerButtonInBuf[9]) && (FM_PS_EN == `PwrSW_Off)) ? 1'b1 : 1'b0;
assign FM_SYS_SIO_PWRBTN_N = PowerButtonOut_ox & PowerbuttonEvtOut;

//----------------------------------------------------------------------
// Internal signal
//----------------------------------------------------------------------
// None

//----------------------------------------------------------------------
// FSM
//----------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Sequential circuit
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Output
//----------------------------------------------------------------------
// None

//----------------------------------------------------------------------
// Internal signal
//----------------------------------------------------------------------
always @ (posedge Strobe125ms or negedge InitResetN) begin
    if(!InitResetN)
        PowerButtonInBuf <= #TD 10'd0;
    else
        PowerButtonInBuf <= #TD {PowerButtonInBuf[8:0], PWR_BTN_IN_N };
end

//----------------------------------------------------------------------
// FSM
//----------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Module instantiation
//--------------------------------------------------------------------------
// None

endmodule // PwrBtnControl
