//******************************************************************************
// File name        : Button.v
// Module name      : Button
// Company          : Caswell
// Project name     : ODS-MR
// Card name        : Yarkon
// Designer         : Fedor Haikin
// Creation Date    : 08.02.2011
// Status           : Under design
// Last modified    : 10.13.2015
// Version          : 1.0
// Description      : This module output debounce button input, interrupt...
// Hierarchy Up     : ODSLS
// Hierarchy Down   :
// Card Release     : 1.0
//******************************************************************************

//------------------------------------------------------------------------------
// Macro define or include file
//------------------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Module declaration
//------------------------------------------------------------------------------
module Button(
    MainReset,      // In, Power or Controller ICH10R Reset
    SlowClock,      // In, Oscillator Clock 32,768 Hz
    Strobe16ms,     // In, Single SlowClock Pulse @ 16 ms
    Strobe125ms,    // In, Single SlowClock Pulse @ 125 ms
    ButtonIn,       // In, Button Input
    Interrupt,      // Out, Single SlowClock Pulse 1s after the button pushed
    StrobeOut,      // Out, Active Wide Strobe 4s after the button pushed
    Release         // Out, Single SlowClock Pulse after the button released
);

//------------------------------------------------------------------------------
// Parameter declaration
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// User defined parameter
//--------------------------------------------------------------------------
parameter RST = 0;

//--------------------------------------------------------------------------
// Standard parameter
//--------------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Local parameter
//--------------------------------------------------------------------------
// time delay, flip-flop output assignment delay for simulation waveform trace
localparam TD = 1;

//------------------------------------------------------------------------------
// Variable declaration
//------------------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Input/Output declaration
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// Input declaration
//--------------------------------------------------------------------------
input           MainReset;
input           SlowClock;
input           Strobe16ms;
input           Strobe125ms;
input           ButtonIn;

//--------------------------------------------------------------------------
// Output declaration
//--------------------------------------------------------------------------
output          Interrupt;
output          Release;
output          StrobeOut;

//------------------------------------------------------------------------------
// Signal declaration
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// Wire declaration
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Combinational, module connection
//----------------------------------------------------------------------
wire            Widest;

//--------------------------------------------------------------------------
// Reg declaration
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Combinational
//----------------------------------------------------------------------
//------------------------------------------------------------------
// Output
//------------------------------------------------------------------
// None

//------------------------------------------------------------------
// Internal signal
//------------------------------------------------------------------
// None

//------------------------------------------------------------------
// FSM
//------------------------------------------------------------------
// None

//----------------------------------------------------------------------
// Sequential
//----------------------------------------------------------------------
//------------------------------------------------------------------
// Output
//------------------------------------------------------------------
reg             Interrupt;
reg             Release;

//------------------------------------------------------------------
// Internal signal
//------------------------------------------------------------------
reg     [2:0]   Debounce; // Debounce shift register
reg             Status;
reg             Strobe;
reg     [5:0]   Timer;

//------------------------------------------------------------------
// FSM
//------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Task/Function description and included task/function description
//------------------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Main code
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// Combinational circuit
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Output
//----------------------------------------------------------------------
assign StrobeOut = RST ? Strobe: Status;

//----------------------------------------------------------------------
// Internal signal
//----------------------------------------------------------------------
assign Widest = Timer[5];

//----------------------------------------------------------------------
// FSM
//----------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Sequential circuit
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Output
//----------------------------------------------------------------------
always @ (posedge SlowClock or negedge MainReset) begin
    if(!MainReset) begin
        Interrupt <= #TD 1'b0;
        Release <= #TD 1'b0;
    end else begin
               Interrupt <= #TD (Timer == 6'h7) & Strobe125ms;
               Release <= #TD (Debounce == 3'h7) & (!Status) & Strobe16ms;
             end
end


//----------------------------------------------------------------------
// Internal signal
//----------------------------------------------------------------------
always @ (posedge SlowClock or negedge MainReset) begin
    if(!MainReset) begin
        Debounce <= #TD 3'h7;
        Status <= #TD 1'b1;
    end else if(Strobe16ms) begin
                  Debounce <= #TD {Debounce[1:0], ButtonIn};
                  Status <= #TD (Debounce == 3'h7) | Status & (Debounce != 3'h0);
              end else begin
                  Debounce <= #TD Debounce;
                  Status <= #TD Status;
              end
end

always @ (posedge SlowClock or negedge MainReset) begin
    if(!MainReset)
        Strobe <= #TD 1'b1;
    else
        Strobe <= #TD (Timer != 6'h1F);
end

always @ (posedge SlowClock or negedge MainReset) begin
    if(!MainReset)
        Timer <= #TD 6'd0;
    else if(Strobe125ms)
           if(Status)
             Timer <= #TD 6'h0;
           else
             Timer <= #TD Widest ? Timer: (Timer + 1'b1);
         else
             Timer <= #TD Timer;
end
//----------------------------------------------------------------------
// FSM
//----------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Module instantiation
//--------------------------------------------------------------------------
// None

endmodule
