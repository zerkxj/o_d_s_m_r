//******************************************************************************
// File name      : LanLED.v
// Module name    : LanLED
// Company        : CASwell
// Project name   : ODS-MR
// Card name      : Ethernet LED
// Designer       : Frank Hsu
// Creation Date  : May 8,2015
// Status         : Under design
// Last modified  : Oct 25,2015
//                :
// Description    : This module controls the Giga Port Speed Leds Colour
// Hierarchy Up   :
// Hierarchy Down :
// Card Release   :
//******************************************************************************

//------------------------------------------------------------------------------
// Macro define or include file
//------------------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Module declaration
//------------------------------------------------------------------------------
module LanLED (
    ALL_PWRGD,  // In, ALL POWER GOOD
    PActivity,  // In, ACT#      signal from LAN controller
    Speed1P,    // In, LINK1000# signal from LAN controller
    Speed2P,    // In, LINK100#  signal from LAN controller
    Speed1R,    // Out, LINK1000# output to BiColor LED
    Speed2R,    // Out, LINK100#  output to BiColor LED
    RActivity   // Out, ACT#      output to LED
);

//------------------------------------------------------------------------------
// Parameter declaration
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// User defined parameter
//--------------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Standard parameter
//--------------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Local parameter
//--------------------------------------------------------------------------
// time delay, flip-flop output assignment delay for simulation waveform trace
localparam TD = 1;

//------------------------------------------------------------------------------
// Variable declaration
//------------------------------------------------------------------------------
integer i_loop;

//------------------------------------------------------------------------------
// Input/Output declaration
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// Input declaration
//--------------------------------------------------------------------------
input           ALL_PWRGD;
input   [1:0]   PActivity;
input   [1:0]   Speed1P;
input   [1:0]   Speed2P;

//--------------------------------------------------------------------------
// Output declaration
//--------------------------------------------------------------------------
output  [1:0]   Speed1R;
output  [1:0]   Speed2R;
output  [1:0]   RActivity;

//------------------------------------------------------------------------------
// Signal declaration
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// Wire declaration
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Combinational, module connection
//----------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Reg declaration
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Combinational
//----------------------------------------------------------------------
//------------------------------------------------------------------
// Output
//------------------------------------------------------------------
reg     [1:0]   RActivity;

//------------------------------------------------------------------
// Internal signal
//------------------------------------------------------------------
// None

//------------------------------------------------------------------
// FSM
//------------------------------------------------------------------
// None

//----------------------------------------------------------------------
// Sequential
//----------------------------------------------------------------------
//------------------------------------------------------------------
// Output
//------------------------------------------------------------------
// None

//------------------------------------------------------------------
// Internal signal
//------------------------------------------------------------------
// None

//------------------------------------------------------------------
// FSM
//------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Task/Function description and included task/function description
//------------------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Main code
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// Combinational circuit
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Output
//----------------------------------------------------------------------
//LinkSpeedLEDs describe the link type of the GigaPhy
//The table below gives the Link modes according to the SpeedLED status
//|Speed1P:Speed2P| LinkMode       |Required LED Color|Speed1R:Speed2R|
//|---------------|----------------|------------------|---------------|
//|        00     | 1000BaseT Link |     Green        |        10     |
//|        01     | 100BaseT Link  |     Orange       |        01     |
//|        10     | 10BaseT Link   |     Orange       |        01     |
//|        11     | NO Link        |     OFF          |        00     |
//|---------------|----------------|------------------|---------------|
assign Speed1R = ALL_PWRGD ? Speed2P: 2'b11;
assign Speed2R = ALL_PWRGD ? Speed1P: 2'b11;

always @ (ALL_PWRGD or Speed1P or Speed2P or PActivity) begin
    for (i_loop=0; i_loop<2; i_loop=i_loop+1) begin
        if (ALL_PWRGD)
            if ({Speed1P[i_loop], Speed2P[i_loop]} == 2'b11)
                RActivity[i_loop] = 1'b1;
            else
                RActivity[i_loop] = ~RActivity[i_loop];
        else
            RActivity[i_loop] = 1'b1;
    end
end

//----------------------------------------------------------------------
// Internal signal
//----------------------------------------------------------------------
// None

//----------------------------------------------------------------------
// FSM
//----------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Sequential circuit
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Output
//----------------------------------------------------------------------
// None

//----------------------------------------------------------------------
// Internal signal
//----------------------------------------------------------------------
// None

//----------------------------------------------------------------------
// FSM
//----------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Module instantiation
//--------------------------------------------------------------------------
// None

endmodule
