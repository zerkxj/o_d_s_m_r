//******************************************************************************
// File name      : InterruptControl.v
// Module name    : InterruptControl
// Company        : Radware
// Project name   : ODS-MR
// Card name      : Yarkon
// Designer       : Fedor Haikin
// Creation Date  : 08.02.2011
// Status         : Under design
// Last modified  : 10.16.2015
// Version        : 1.0
// Description    : This module controls Interrupts
// Hierarchy Up   : ODS_MR
// Hierarchy Down : ---
// Card Release   : 1.0
//******************************************************************************
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Macro define or include file
//------------------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Module declaration
//------------------------------------------------------------------------------
module InterruptControl (
    WatchDogIREQ,       // In, Watch Dog Interrupt Request
    Wr,                 // In, LPC write signal
    Addr,               // In, LPC register address
    DataIntReg,         // In, Interrupt register(0x09)
    DataWr,             // In, Data to be written to register
    Interrupt,          // In, Power & Reset Interrupts and Button release
    InterruptRegister,  // Out, Interrupt Control / Status Register
    InterruptD          // Out, Interrupt Request to CPU
);

//------------------------------------------------------------------------------
// Parameter declaration
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// User defined parameter
//--------------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Standard parameter
//--------------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Local parameter
//--------------------------------------------------------------------------
// time delay, flip-flop output assignment delay for simulation waveform trace
localparam TD = 1;

//------------------------------------------------------------------------------
// Variable declaration
//------------------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Input/Output declaration
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// Input declaration
//--------------------------------------------------------------------------
input           WatchDogIREQ;
input           Wr;
input   [7:0]   Addr;
input   [7:0]   DataIntReg;
input   [7:0]   DataWr;
input   [3:0]   Interrupt;

//--------------------------------------------------------------------------
// Output declaration
//--------------------------------------------------------------------------
output  [6:4]   InterruptRegister;
output          InterruptD;

//------------------------------------------------------------------------------
// Signal declaration
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// Wire declaration
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Combinational, module connection
//----------------------------------------------------------------------
wire            ATX;
wire    [2:0]   EnableInt;
wire            ResetEvent;
wire            PowerEvent;
wire            WrRegInt;
wire    [6:4]   ClearInterrupt;
wire            IREQWatchDog;
wire            IREQResetButton;
wire            IREQPwrButton;
wire            InterruptRequest;

//--------------------------------------------------------------------------
// Reg declaration
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Combinational
//----------------------------------------------------------------------
//------------------------------------------------------------------
// Output
//------------------------------------------------------------------
// None

//------------------------------------------------------------------
// Internal signal
//------------------------------------------------------------------
// None

//------------------------------------------------------------------
// FSM
//------------------------------------------------------------------
// None

//----------------------------------------------------------------------
// Sequential
//----------------------------------------------------------------------
//------------------------------------------------------------------
// Output
//------------------------------------------------------------------
// None

//------------------------------------------------------------------
// Internal signal
//------------------------------------------------------------------
// None

//------------------------------------------------------------------
// FSM
//------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Task/Function description and included task/function description
//------------------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Main code
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// Combinational circuit
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Output
//----------------------------------------------------------------------
assign InterruptRegister = {IREQWatchDog, IREQResetButton, IREQPwrButton};

assign InterruptD = InterruptRequest ? 1'b0 : 1'bz;


//----------------------------------------------------------------------
// Internal signal
//----------------------------------------------------------------------
assign ATX = DataIntReg[3];
assign EnableInt = DataIntReg[2:0];
assign ResetEvent = ATX ? Interrupt[0] : Interrupt[1];
assign PowerEvent = ATX ? Interrupt[2] : Interrupt[3];
assign WrRegInt = Wr & (Addr == 8'h09);
assign ClearInterrupt = DataWr[6:4] & {3{WrRegInt}};
assign IREQWatchDog = WatchDogIREQ | DataIntReg[6];
assign IREQResetButton = ResetEvent | DataIntReg[5] & (!ClearInterrupt[5]);
assign IREQPwrButton = PowerEvent | DataIntReg[4] & (!ClearInterrupt[4]);
assign InterruptRequest = |({IREQWatchDog, IREQResetButton, IREQPwrButton} &
                            EnableInt);

//----------------------------------------------------------------------
// FSM
//----------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Sequential circuit
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Output
//----------------------------------------------------------------------
// None

//----------------------------------------------------------------------
// Internal signal
//----------------------------------------------------------------------
// None

//----------------------------------------------------------------------
// FSM
//----------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Module instantiation
//--------------------------------------------------------------------------
// None

endmodule
