///////////////////////////////////////////////////////////////////
// File name      : OpenDrain.v
// Module name    : OpenDrain
// Company        : Radware
// Project name   : Mekong XGE
// Card name      : MMBXGE
// Designer       : Fedor Haikin
// Creation Date  : 08.05.2007
// Status         : Under design
// Last modified  : 25.06.2007
// Altera Version : 1.0
// Description    : This module provides individual bus signal Open Drain Control
// Hierarchy Up	  : MuxDisplay
// Hierarchy Down : ---
// Card Release	  : 1.0
///////////////////////////////////////////////////////////////////
`ifdef		OpenDrain
`else
`define		OpenDrain
///////////////////////////////////////////////////////////////////
module	OpenDrain(
	Control,			// Output Buffer Control
	DataOut
	);
///////////////////////////////////////////////////////////////////
parameter	Width = 8;
///////////////////////////////////////////////////////////////////
input	[Width:1]	Control;
output	[Width:1]	DataOut;
///////////////////////////////////////////////////////////////////
reg		[Width:1]	DataOut;
integer				Loop;
///////////////////////////////////////////////////////////////////
always	@(Control)
  for(Loop = 1; Loop <= Width; Loop = Loop + 1)
     //DataOut[Loop] = Control[Loop] ? 1'b0 : 1'bz;
     DataOut[Loop] = Control[Loop] ? 1'b0 : 1'b1;
///////////////////////////////////////////////////////////////////
endmodule
///////////////////////////////////////////////////////////////////
`endif
