//******************************************************************************
// File name      : FanDisplay.v
// Module name    : FanDisplay
// Company        : Radware
// Project name   : ODS-MR
// Card name      : Yarkon
// Designer       : Fedor Haikin
// Creation Date  : 12.04.2011
// Status         : Under design
// Last modified  : 10.26.2015
// Version        : 1.0
// Description    : This module controls FAN Status LED
// Hierarchy Up   : ODS_MR
// Hierarchy Down : -------
// Card Release   : 1.0
//******************************************************************************

//------------------------------------------------------------------------------
// Macro define or include file
//------------------------------------------------------------------------------
`define FANLedOff 2'b11
`define FANLedRed 2'b10
`define FANLedGreen 2'b01

//------------------------------------------------------------------------------
// Module declaration
//------------------------------------------------------------------------------
module FanLED (
    SlowClock,      // In, Oscillator Clock 32,768 Hz
    Reset_N,        // In, reset
    Strobe16ms,     // In, Single SlowClock Pulse @ 16 ms
    Beep,           // In, Fan Fail - 1, FanOK - 0; - has internal weak P/U
    FanLedCtrlReg,  // In, Fan LED control register

    FanFail,        // Out, Fan Led indication
    FanOK           // Out, Fan Led indication
);

//------------------------------------------------------------------------------
// Parameter declaration
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// User defined parameter
//--------------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Standard parameter
//--------------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Local parameter
//--------------------------------------------------------------------------
// time delay, flip-flop output assignment delay for simulation waveform trace
localparam TD = 1;

//------------------------------------------------------------------------------
// Variable declaration
//------------------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Input/Output declaration
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// Input declaration
//--------------------------------------------------------------------------
input           SlowClock;
input           Reset_N;
input           Strobe16ms;
input           Beep;
input   [3:0]   FanLedCtrlReg;

//--------------------------------------------------------------------------
// Output declaration
//--------------------------------------------------------------------------
output          FanFail;
output          FanOK;

//------------------------------------------------------------------------------
// Signal declaration
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// Wire declaration
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Combinational, module connection
//----------------------------------------------------------------------
wire            Fail;

//--------------------------------------------------------------------------
// Reg declaration
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Combinational
//----------------------------------------------------------------------
//------------------------------------------------------------------
// Output
//------------------------------------------------------------------
reg             FanFail;
reg             FanOK;

//------------------------------------------------------------------
// Internal signal
//------------------------------------------------------------------
reg             Tone;
reg     [1:0]   Sample;
reg             FanFailx;
reg             FanOKx;

//------------------------------------------------------------------
// FSM
//------------------------------------------------------------------
// None

//----------------------------------------------------------------------
// Sequential
//----------------------------------------------------------------------
//------------------------------------------------------------------
// Output
//------------------------------------------------------------------
// None

//------------------------------------------------------------------
// Internal signal
//------------------------------------------------------------------
// None

//------------------------------------------------------------------
// FSM
//------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Task/Function description and included task/function description
//------------------------------------------------------------------------------
// None

//------------------------------------------------------------------------------
// Main code
//------------------------------------------------------------------------------
//--------------------------------------------------------------------------
// Combinational circuit
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Output
//----------------------------------------------------------------------
always @ (FanLedCtrlReg or FanOKx or FanFailx) begin
    casex (FanLedCtrlReg)
        4'bxxx0: {FanOK, FanFail} = {FanOKx, FanFailx};
        4'bxx11: {FanOK, FanFail} = `FANLedOff;
        4'bx111: {FanOK, FanFail} = `FANLedGreen;
        4'b1111: {FanOK, FanFail} = `FANLedRed;
        default: {FanOK, FanFail} = `FANLedOff;
    endcase
end

//----------------------------------------------------------------------
// Internal signal
//----------------------------------------------------------------------
assign Fail = |Sample;

//----------------------------------------------------------------------
// FSM
//----------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Sequential circuit
//--------------------------------------------------------------------------
//----------------------------------------------------------------------
// Output
//----------------------------------------------------------------------
// None

//----------------------------------------------------------------------
// Internal signal
//----------------------------------------------------------------------
always @ (negedge Reset_N or posedge SlowClock) begin
    if (!Reset_N)
        Sample <= #TD 2'd0;
    else if (Tone)
             Sample <= #TD 2'd3;
         else if (Strobe16ms & Fail)
                  Sample <= #TD Sample - 2'd1;
              else
                  Sample <= #TD Sample;
end

always @ (negedge Reset_N or posedge SlowClock) begin
    if (!Reset_N) begin
        Tone <= #TD 1'b0;
        FanFailx <= #TD 1'b0;
        FanOKx <= #TD 1'b0;
    end else begin
        Tone <= #TD Beep;
        FanFailx <= #TD Fail;
        FanOKx <= #TD !Fail;
    end
end

//----------------------------------------------------------------------
// FSM
//----------------------------------------------------------------------
// None

//--------------------------------------------------------------------------
// Module instantiation
//--------------------------------------------------------------------------
// None

endmodule
